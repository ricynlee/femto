    assign array[0] = 32'h10001197;
    assign array[1] = 32'h80018193;
    assign array[2] = 32'h10000117;
    assign array[3] = 32'h1f810113;
    assign array[4] = 32'h11712009;
    assign array[5] = 32'h0040c022;
    assign array[6] = 32'hf00007b7;
    assign array[7] = 32'h00078023;
    assign array[8] = 32'h0000a001;
    assign array[9] = 32'h00000014;
    assign array[10] = 32'h00000000;
    assign array[11] = 32'h00527a01;
    assign array[12] = 32'h01017c01;
    assign array[13] = 32'h07020d1b;
    assign array[14] = 32'h00000001;
    assign array[15] = 32'h00000010;
    assign array[16] = 32'h0000001c;
    assign array[17] = 32'hffffffbc;
    assign array[18] = 32'h00000012;
    assign array[19] = 32'h00000000;
