
module dbusif (
    input clk,
    input rstn,

);

endmodule
