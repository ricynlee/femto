    assign array[0] = 32'h10004117;
    assign array[1] = 32'h00010113;
    assign array[2] = 32'h06a0006f;
    assign array[3] = 32'hc2221151;
    assign array[4] = 32'h440dc406;
    assign array[5] = 32'h45854601;
    assign array[6] = 32'h2a9d4501;
    assign array[7] = 32'h00040537;
    assign array[8] = 32'h46012285;
    assign array[9] = 32'h45014581;
    assign array[10] = 32'h053722a5;
    assign array[11] = 32'h147d0004;
    assign array[12] = 32'hf06d2a81;
    assign array[13] = 32'h441240a2;
    assign array[14] = 32'h80820131;
    assign array[15] = 32'hc2221151;
    assign array[16] = 32'hc026c406;
    assign array[17] = 32'h10000437;
    assign array[18] = 32'he91920dd;
    assign array[19] = 32'hfd6d2235;
    assign array[20] = 32'h44123f75;
    assign array[21] = 32'h448240a2;
    assign array[22] = 32'h10000337;
    assign array[23] = 32'h83020131;
    assign array[24] = 32'h20d58522;
    assign array[25] = 32'h00140493;
    assign array[26] = 32'h00080537;
    assign array[27] = 32'h84262211;
    assign array[28] = 32'h1141bfe1;
    assign array[29] = 32'hc422c606;
    assign array[30] = 32'h2281c226;
    assign array[31] = 32'h4481287d;
    assign array[32] = 32'ha81dc002;
    assign array[33] = 32'h10000513;
    assign array[34] = 32'h20fd20e5;
    assign array[35] = 32'h4782e905;
    assign array[36] = 32'h0087a7b3;
    assign array[37] = 32'h0017c593;
    assign array[38] = 32'hf593c099;
    assign array[39] = 32'h46010ff7;
    assign array[40] = 32'h20fd4501;
    assign array[41] = 32'h07930405;
    assign array[42] = 32'h1de30400;
    assign array[43] = 32'h4782fcf4;
    assign array[44] = 32'hc03e0785;
    assign array[45] = 32'h00878e63;
    assign array[46] = 32'hb7e94401;
    assign array[47] = 32'hd571288d;
    assign array[48] = 32'h287d4521;
    assign array[49] = 32'h45814601;
    assign array[50] = 32'h20d94501;
    assign array[51] = 32'ha0013f85;
    assign array[52] = 32'hf4d5e481;
    assign array[53] = 32'hb76d4485;
    assign array[54] = 32'h00030537;
    assign array[55] = 32'h28692851;
    assign array[56] = 32'h20b1d96d;
    assign array[57] = 32'hbfe9dd6d;
    assign array[58] = 32'h400007b7;
    assign array[59] = 32'h470543dc;
    assign array[60] = 32'h00a71533;
    assign array[61] = 32'h00e59763;
    assign array[62] = 32'h07378fc9;
    assign array[63] = 32'hc35c4000;
    assign array[64] = 32'h45138082;
    assign array[65] = 32'h8fe9fff5;
    assign array[66] = 32'h4785bfcd;
    assign array[67] = 32'h00a79533;
    assign array[68] = 32'h0737c599;
    assign array[69] = 32'h431c4000;
    assign array[70] = 32'hc3088d5d;
    assign array[71] = 32'h07b78082;
    assign array[72] = 32'h43984000;
    assign array[73] = 32'hfff54513;
    assign array[74] = 32'hc3888d79;
    assign array[75] = 32'h07b78082;
    assign array[76] = 32'hc5035000;
    assign array[77] = 32'h89050037;
    assign array[78] = 32'h07b78082;
    assign array[79] = 32'h47095000;
    assign array[80] = 32'h00e781a3;
    assign array[81] = 32'he9018082;
    assign array[82] = 32'h80824501;
    assign array[83] = 32'h40a24501;
    assign array[84] = 32'h01314412;
    assign array[85] = 32'h11518082;
    assign array[86] = 32'hc406c222;
    assign array[87] = 32'h3fc1842a;
    assign array[88] = 32'h07b7d575;
    assign array[89] = 32'hc7835000;
    assign array[90] = 32'h00230017;
    assign array[91] = 32'hb7c500f4;
    assign array[92] = 32'h700007b7;
    assign array[93] = 32'h8082c388;
    assign array[94] = 32'h700007b7;
    assign array[95] = 32'h80824388;
    assign array[96] = 32'h700007b7;
    assign array[97] = 32'h0737c388;
    assign array[98] = 32'h431c7000;
    assign array[99] = 32'h8082fffd;
    assign array[100] = 32'hc4221141;
    assign array[101] = 32'h4593842e;
    assign array[102] = 32'h45050015;
    assign array[103] = 32'hc032c606;
    assign array[104] = 32'h459337ad;
    assign array[105] = 32'h45090014;
    assign array[106] = 32'h4602378d;
    assign array[107] = 32'h40b24422;
    assign array[108] = 32'h00164593;
    assign array[109] = 32'h0141450d;
    assign array[110] = 32'h1151bf89;
    assign array[111] = 32'h45814601;
    assign array[112] = 32'hc4064501;
    assign array[113] = 32'h458137f1;
    assign array[114] = 32'h3f394501;
    assign array[115] = 32'h45054585;
    assign array[116] = 32'h45853f21;
    assign array[117] = 32'h3f094509;
    assign array[118] = 32'h458540a2;
    assign array[119] = 32'h0131450d;
    assign array[120] = 32'h0000b721;
