    assign array[0] = 32'h10001197;
    assign array[1] = 32'h80018193;
    assign array[2] = 32'h10000117;
    assign array[3] = 32'h1f810113;
    assign array[4] = 32'h28812019;
    assign array[5] = 32'h11412855;
    assign array[6] = 32'h0800c622;
    assign array[7] = 32'h00000793;
    assign array[8] = 32'hfef42a23;
    assign array[9] = 32'h100007b7;
    assign array[10] = 32'h00078793;
    assign array[11] = 32'hfef42823;
    assign array[12] = 32'hfe042c23;
    assign array[13] = 32'h2703a829;
    assign array[14] = 32'h2783ff04;
    assign array[15] = 32'h97baff84;
    assign array[16] = 32'h00078023;
    assign array[17] = 32'hff842783;
    assign array[18] = 32'h2c230785;
    assign array[19] = 32'h2703fef4;
    assign array[20] = 32'h2783ff84;
    assign array[21] = 32'h60e3ff44;
    assign array[22] = 32'h0001fef7;
    assign array[23] = 32'h01414432;
    assign array[24] = 32'h11318082;
    assign array[25] = 32'h0840c822;
    assign array[26] = 32'h00000793;
    assign array[27] = 32'hfef42a23;
    assign array[28] = 32'h1ec00793;
    assign array[29] = 32'hfef42823;
    assign array[30] = 32'h100007b7;
    assign array[31] = 32'h00078793;
    assign array[32] = 32'hfef42623;
    assign array[33] = 32'hfe042c23;
    assign array[34] = 32'h2703a035;
    assign array[35] = 32'h2783ff04;
    assign array[36] = 32'h973eff84;
    assign array[37] = 32'hfec42683;
    assign array[38] = 32'hff842783;
    assign array[39] = 32'h470397b6;
    assign array[40] = 32'h77130007;
    assign array[41] = 32'h80230ff7;
    assign array[42] = 32'h278300e7;
    assign array[43] = 32'h0785ff84;
    assign array[44] = 32'hfef42c23;
    assign array[45] = 32'hff842703;
    assign array[46] = 32'hff442783;
    assign array[47] = 32'hfcf767e3;
    assign array[48] = 32'h44420001;
    assign array[49] = 32'h80820151;
    assign array[50] = 32'hcc061111;
    assign array[51] = 32'h0860ca22;
    assign array[52] = 32'h400007b7;
    assign array[53] = 32'hc3d84709;
    assign array[54] = 32'h400007b7;
    assign array[55] = 32'hc3984709;
    assign array[56] = 32'hfe042823;
    assign array[57] = 32'h2783a031;
    assign array[58] = 32'h0785ff04;
    assign array[59] = 32'hfef42823;
    assign array[60] = 32'hff042703;
    assign array[61] = 32'h879367e1;
    assign array[62] = 32'hc96369f7;
    assign array[63] = 32'h07b700e7;
    assign array[64] = 32'hc7835000;
    assign array[65] = 32'hf7930037;
    assign array[66] = 32'hfff10ff7;
    assign array[67] = 32'h500007b7;
    assign array[68] = 32'h0037c783;
    assign array[69] = 32'h0ff7f793;
    assign array[70] = 32'h07b7cb89;
    assign array[71] = 32'h43984000;
    assign array[72] = 32'h400007b7;
    assign array[73] = 32'h00274713;
    assign array[74] = 32'h07b7c398;
    assign array[75] = 32'hc7835000;
    assign array[76] = 32'hf7930037;
    assign array[77] = 32'hf7cd0ff7;
    assign array[78] = 32'h400007b7;
    assign array[79] = 32'h0007a023;
    assign array[80] = 32'h400007b7;
    assign array[81] = 32'h0007a223;
    assign array[82] = 32'h200007b7;
    assign array[83] = 32'hfef42623;
    assign array[84] = 32'h50000737;
    assign array[85] = 32'hfec42783;
    assign array[86] = 32'h00178693;
    assign array[87] = 32'hfed42623;
    assign array[88] = 32'h00174703;
    assign array[89] = 32'h0ff77713;
    assign array[90] = 32'h00e78023;
    assign array[91] = 32'hfe042423;
    assign array[92] = 32'h2783a031;
    assign array[93] = 32'h0785fe84;
    assign array[94] = 32'hfef42423;
    assign array[95] = 32'hfe842703;
    assign array[96] = 32'h000f47b7;
    assign array[97] = 32'h23f78793;
    assign array[98] = 32'h00e7c963;
    assign array[99] = 32'h500007b7;
    assign array[100] = 32'h0037c783;
    assign array[101] = 32'h0ff7f793;
    assign array[102] = 32'h07b7ffe9;
    assign array[103] = 32'hc7835000;
    assign array[104] = 32'hf7930037;
    assign array[105] = 32'hd7cd0ff7;
    assign array[106] = 32'h200007b7;
    assign array[107] = 32'hfef42223;
    assign array[108] = 32'hfe442783;
    assign array[109] = 32'ha0019782;
    assign array[110] = 32'h00000014;
    assign array[111] = 32'h00000000;
    assign array[112] = 32'h00527a01;
    assign array[113] = 32'h01017c01;
    assign array[114] = 32'h07020d1b;
    assign array[115] = 32'h00000001;
    assign array[116] = 32'h00000010;
    assign array[117] = 32'h0000001c;
    assign array[118] = 32'hfffffe28;
    assign array[119] = 32'h00000016;
    assign array[120] = 32'h00000000;
    assign array[121] = 32'h40000000;
    assign array[122] = 32'h50000000;
