module wrapper();
    // clk_gen clk_gen
    // (
    //     .clk_out(clk),
    //     .clk_in(sysclk)
    // );
    
endmodule
