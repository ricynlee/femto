module ioring();

endmodule
