    assign array[0] = 32'h10001197;
    assign array[1] = 32'h80018193;
    assign array[2] = 32'h10000117;
    assign array[3] = 32'h1f810113;
    assign array[4] = 32'h117120e9;
    assign array[5] = 32'h0040c022;
    assign array[6] = 32'h700007b7;
    assign array[7] = 32'h50415737;
    assign array[8] = 32'h35370713;
    assign array[9] = 32'ha001c398;
    assign array[10] = 32'hc0221171;
    assign array[11] = 32'h07b70040;
    assign array[12] = 32'h57377000;
    assign array[13] = 32'h07134641;
    assign array[14] = 32'hc39894c7;
    assign array[15] = 32'h1161a001;
    assign array[16] = 32'h0020c222;
    assign array[17] = 32'hfea42c23;
    assign array[18] = 32'h700007b7;
    assign array[19] = 32'hff842703;
    assign array[20] = 32'h0001c398;
    assign array[21] = 32'h01214412;
    assign array[22] = 32'h11618082;
    assign array[23] = 32'h0020c222;
    assign array[24] = 32'h0da387aa;
    assign array[25] = 32'h4703fef4;
    assign array[26] = 32'h57b7ffb4;
    assign array[27] = 32'h87935052;
    assign array[28] = 32'h8f5de007;
    assign array[29] = 32'h700007b7;
    assign array[30] = 32'h0001c398;
    assign array[31] = 32'h01214412;
    assign array[32] = 32'h11518082;
    assign array[33] = 32'h0060c422;
    assign array[34] = 32'hfea42a23;
    assign array[35] = 32'hff442783;
    assign array[36] = 32'hfef42c23;
    assign array[37] = 32'h2783a01d;
    assign array[38] = 32'hc783ff84;
    assign array[39] = 32'h873e0007;
    assign array[40] = 32'h505257b7;
    assign array[41] = 32'he0078793;
    assign array[42] = 32'h07b78f5d;
    assign array[43] = 32'hc3987000;
    assign array[44] = 32'hff842783;
    assign array[45] = 32'h2c230785;
    assign array[46] = 32'h2783fef4;
    assign array[47] = 32'hc783ff84;
    assign array[48] = 32'hfbf10007;
    assign array[49] = 32'h700007b7;
    assign array[50] = 32'h50525737;
    assign array[51] = 32'he0a70713;
    assign array[52] = 32'h0001c398;
    assign array[53] = 32'h01314422;
    assign array[54] = 32'h11518082;
    assign array[55] = 32'hc222c406;
    assign array[56] = 32'h07b70060;
    assign array[57] = 32'h47052000;
    assign array[58] = 32'h00e78023;
    assign array[59] = 32'h700007b7;
    assign array[60] = 32'hc3984719;
    assign array[61] = 32'h700007b7;
    assign array[62] = 32'h08000713;
    assign array[63] = 32'h4505c3d8;
    assign array[64] = 32'h000120a9;
    assign array[65] = 32'h200007b7;
    assign array[66] = 32'h0007c783;
    assign array[67] = 32'h3711ffe5;
    assign array[68] = 32'h40a20001;
    assign array[69] = 32'h01314412;
    assign array[70] = 32'h11718082;
    assign array[71] = 32'h0040c022;
    assign array[72] = 32'h200007b7;
    assign array[73] = 32'h00078023;
    assign array[74] = 32'h44020001;
    assign array[75] = 32'h80820111;
    assign array[76] = 32'hc2221161;
    assign array[77] = 32'h2c230020;
    assign array[78] = 32'h2783fea4;
    assign array[79] = 32'h9073ff84;
    assign array[80] = 32'h00013057;
    assign array[81] = 32'h01214412;
    assign array[82] = 32'h11418082;
    assign array[83] = 32'hc422c606;
    assign array[84] = 32'h87aa0800;
    assign array[85] = 32'hfef409a3;
    assign array[86] = 32'hff344783;
    assign array[87] = 32'h0513c799;
    assign array[88] = 32'h37f91780;
    assign array[89] = 32'h30046073;
    assign array[90] = 32'h7073a019;
    assign array[91] = 32'h00013004;
    assign array[92] = 32'h442240b2;
    assign array[93] = 32'h80820141;
    assign array[94] = 32'hfd410113;
    assign array[95] = 32'hd216d406;
    assign array[96] = 32'hce1ed01a;
    assign array[97] = 32'hca2acc22;
    assign array[98] = 32'hc632c82e;
    assign array[99] = 32'hc23ac436;
    assign array[100] = 32'h1060c03e;
    assign array[101] = 32'h00013759;
    assign array[102] = 32'h529250a2;
    assign array[103] = 32'h43f25302;
    assign array[104] = 32'h45524462;
    assign array[105] = 32'h463245c2;
    assign array[106] = 32'h471246a2;
    assign array[107] = 32'h01134782;
    assign array[108] = 32'h007302c1;
    assign array[109] = 32'h00003020;
    assign array[110] = 32'h00000014;
    assign array[111] = 32'h00000000;
    assign array[112] = 32'h00527a01;
    assign array[113] = 32'h01017c01;
    assign array[114] = 32'h07020d1b;
    assign array[115] = 32'h00000001;
    assign array[116] = 32'h00000010;
    assign array[117] = 32'h0000001c;
    assign array[118] = 32'hfffffe28;
    assign array[119] = 32'h00000012;
    assign array[120] = 32'h00000000;
