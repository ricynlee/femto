`ifndef TIMESCALE_HEADER
`define TIMESCALE_HEADER

`timescale 1ns/1ps

`endif // TIMESCALE_HEADER
