    assign array[0] = 32'h10001197;
    assign array[1] = 32'h80018193;
    assign array[2] = 32'h10000117;
    assign array[3] = 32'h1f810113;
    assign array[4] = 32'h159000ef;
    assign array[5] = 32'h600007b7;
    assign array[6] = 32'h30000713;
    assign array[7] = 32'h00e79323;
    assign array[8] = 32'h03374609;
    assign array[9] = 32'h22833000;
    assign array[10] = 32'h82230003;
    assign array[11] = 32'h82a300c7;
    assign array[12] = 32'h450d00c7;
    assign array[13] = 32'h00a78123;
    assign array[14] = 32'h00078123;
    assign array[15] = 32'h00078123;
    assign array[16] = 32'h00078123;
    assign array[17] = 32'h11100593;
    assign array[18] = 32'h00b79023;
    assign array[19] = 32'h90234745;
    assign array[20] = 32'h470500e7;
    assign array[21] = 32'h00e79023;
    assign array[22] = 32'h00079023;
    assign array[23] = 32'h0037c383;
    assign array[24] = 32'h0037c683;
    assign array[25] = 32'h0037c703;
    assign array[26] = 32'h06e203c2;
    assign array[27] = 32'h00d3e3b3;
    assign array[28] = 32'h0037c683;
    assign array[29] = 32'h0083d393;
    assign array[30] = 32'h67330762;
    assign array[31] = 32'h83210077;
    assign array[32] = 32'h82a306e2;
    assign array[33] = 32'h8f5500c7;
    assign array[34] = 32'h00e28a63;
    assign array[35] = 32'h464157b7;
    assign array[36] = 32'h70000737;
    assign array[37] = 32'h94c78793;
    assign array[38] = 32'ha001c31c;
    assign array[39] = 32'h00435683;
    assign array[40] = 32'h00c78223;
    assign array[41] = 32'h00a78123;
    assign array[42] = 32'h00b79023;
    assign array[43] = 32'h600007b7;
    assign array[44] = 32'h0007d703;
    assign array[45] = 32'hff6d8b09;
    assign array[46] = 32'h00078123;
    assign array[47] = 32'h00078123;
    assign array[48] = 32'h81234711;
    assign array[49] = 32'h474500e7;
    assign array[50] = 32'h00e79023;
    assign array[51] = 32'h600007b7;
    assign array[52] = 32'h0007d703;
    assign array[53] = 32'hff6d8b09;
    assign array[54] = 32'h82a34709;
    assign array[55] = 32'h470500e7;
    assign array[56] = 32'h00e79023;
    assign array[57] = 32'h60000737;
    assign array[58] = 32'h00075783;
    assign array[59] = 32'hffed8b89;
    assign array[60] = 32'h00071023;
    assign array[61] = 32'h00374603;
    assign array[62] = 32'h00374783;
    assign array[63] = 32'h02a34589;
    assign array[64] = 32'h07a200b7;
    assign array[65] = 32'h8a638fd1;
    assign array[66] = 32'h57b700f6;
    assign array[67] = 32'h07374641;
    assign array[68] = 32'h87937000;
    assign array[69] = 32'hc31c94c7;
    assign array[70] = 32'h8082a001;
    assign array[71] = 32'h07b76705;
    assign array[72] = 32'h06936000;
    assign array[73] = 32'h9323b807;
    assign array[74] = 32'h460900d7;
    assign array[75] = 32'h30000337;
    assign array[76] = 32'h00032283;
    assign array[77] = 32'h00c78223;
    assign array[78] = 32'h00c782a3;
    assign array[79] = 32'h8123452d;
    assign array[80] = 32'h812300a7;
    assign array[81] = 32'h81230007;
    assign array[82] = 32'h81230007;
    assign array[83] = 32'h05930007;
    assign array[84] = 32'h90231110;
    assign array[85] = 32'h46c500b7;
    assign array[86] = 32'h00d79023;
    assign array[87] = 32'h82170713;
    assign array[88] = 32'h00e79023;
    assign array[89] = 32'h90234705;
    assign array[90] = 32'h902300e7;
    assign array[91] = 32'hc3830007;
    assign array[92] = 32'hc6830037;
    assign array[93] = 32'hc7030037;
    assign array[94] = 32'h03c20037;
    assign array[95] = 32'he3b306e2;
    assign array[96] = 32'hc68300d3;
    assign array[97] = 32'hd3930037;
    assign array[98] = 32'h07620083;
    assign array[99] = 32'h00776733;
    assign array[100] = 32'h06e28321;
    assign array[101] = 32'h00c782a3;
    assign array[102] = 32'h8a638f55;
    assign array[103] = 32'h57b700e2;
    assign array[104] = 32'h07374641;
    assign array[105] = 32'h87937000;
    assign array[106] = 32'hc31c94c7;
    assign array[107] = 32'h5683a001;
    assign array[108] = 32'h82230043;
    assign array[109] = 32'h812300c7;
    assign array[110] = 32'h902300a7;
    assign array[111] = 32'h07b700b7;
    assign array[112] = 32'hd7036000;
    assign array[113] = 32'h8b090007;
    assign array[114] = 32'h8123ff6d;
    assign array[115] = 32'h81230007;
    assign array[116] = 32'h47110007;
    assign array[117] = 32'h00e78123;
    assign array[118] = 32'h90234745;
    assign array[119] = 32'h073700e7;
    assign array[120] = 32'h57836000;
    assign array[121] = 32'h8b890007;
    assign array[122] = 32'h6785ffed;
    assign array[123] = 32'h82178793;
    assign array[124] = 32'h00f71023;
    assign array[125] = 32'h600007b7;
    assign array[126] = 32'h0007d703;
    assign array[127] = 32'hff6d8b09;
    assign array[128] = 32'h82a34709;
    assign array[129] = 32'h470500e7;
    assign array[130] = 32'h00e79023;
    assign array[131] = 32'h60000737;
    assign array[132] = 32'h00075783;
    assign array[133] = 32'hffed8b89;
    assign array[134] = 32'h00071023;
    assign array[135] = 32'h00374603;
    assign array[136] = 32'h00374783;
    assign array[137] = 32'h02a34589;
    assign array[138] = 32'h07a200b7;
    assign array[139] = 32'h8a638fd1;
    assign array[140] = 32'h57b700f6;
    assign array[141] = 32'h07374641;
    assign array[142] = 32'h87937000;
    assign array[143] = 32'hc31c94c7;
    assign array[144] = 32'h8082a001;
    assign array[145] = 32'h07b76711;
    assign array[146] = 32'h07136000;
    assign array[147] = 32'h9323b817;
    assign array[148] = 32'h460900e7;
    assign array[149] = 32'h30000337;
    assign array[150] = 32'h00032283;
    assign array[151] = 32'h00c78223;
    assign array[152] = 32'h00c782a3;
    assign array[153] = 32'h03b00513;
    assign array[154] = 32'h00a78123;
    assign array[155] = 32'h00078123;
    assign array[156] = 32'h00078123;
    assign array[157] = 32'h00078123;
    assign array[158] = 32'h11100593;
    assign array[159] = 32'h00b79023;
    assign array[160] = 32'h90234745;
    assign array[161] = 32'h670500e7;
    assign array[162] = 32'h82170713;
    assign array[163] = 32'h00e79023;
    assign array[164] = 32'h04100713;
    assign array[165] = 32'h00e79023;
    assign array[166] = 32'h00079023;
    assign array[167] = 32'h0037c383;
    assign array[168] = 32'h0037c683;
    assign array[169] = 32'h0037c703;
    assign array[170] = 32'h06e203c2;
    assign array[171] = 32'h00d3e3b3;
    assign array[172] = 32'h0037c683;
    assign array[173] = 32'h0083d393;
    assign array[174] = 32'h67330762;
    assign array[175] = 32'h83210077;
    assign array[176] = 32'h82a306e2;
    assign array[177] = 32'h8f5500c7;
    assign array[178] = 32'h00e28a63;
    assign array[179] = 32'h464157b7;
    assign array[180] = 32'h70000737;
    assign array[181] = 32'h94c78793;
    assign array[182] = 32'ha001c31c;
    assign array[183] = 32'h00435683;
    assign array[184] = 32'h00c78223;
    assign array[185] = 32'h00a78123;
    assign array[186] = 32'h00b79023;
    assign array[187] = 32'h600007b7;
    assign array[188] = 32'h0007d703;
    assign array[189] = 32'hff6d8b09;
    assign array[190] = 32'h00078123;
    assign array[191] = 32'h00078123;
    assign array[192] = 32'h81234711;
    assign array[193] = 32'h474500e7;
    assign array[194] = 32'h00e79023;
    assign array[195] = 32'h60000737;
    assign array[196] = 32'h00075783;
    assign array[197] = 32'hffed8b89;
    assign array[198] = 32'h87936785;
    assign array[199] = 32'h10238217;
    assign array[200] = 32'h07b700f7;
    assign array[201] = 32'hd7036000;
    assign array[202] = 32'h8b090007;
    assign array[203] = 32'h4709ff6d;
    assign array[204] = 32'h00e782a3;
    assign array[205] = 32'h04100713;
    assign array[206] = 32'h00e79023;
    assign array[207] = 32'h60000737;
    assign array[208] = 32'h00075783;
    assign array[209] = 32'hffed8b89;
    assign array[210] = 32'h00071023;
    assign array[211] = 32'h00374603;
    assign array[212] = 32'h00374783;
    assign array[213] = 32'h02a34589;
    assign array[214] = 32'h07a200b7;
    assign array[215] = 32'h8a638fd1;
    assign array[216] = 32'h57b700f6;
    assign array[217] = 32'h07374641;
    assign array[218] = 32'h87937000;
    assign array[219] = 32'hc31c94c7;
    assign array[220] = 32'h8082a001;
    assign array[221] = 32'h07b77771;
    assign array[222] = 32'h07136000;
    assign array[223] = 32'h9323b437;
    assign array[224] = 32'h460900e7;
    assign array[225] = 32'h30000337;
    assign array[226] = 32'h00032283;
    assign array[227] = 32'h00c78223;
    assign array[228] = 32'h00c782a3;
    assign array[229] = 32'hfbb00513;
    assign array[230] = 32'h00a78123;
    assign array[231] = 32'h00078123;
    assign array[232] = 32'h00078123;
    assign array[233] = 32'h00078123;
    assign array[234] = 32'h11100593;
    assign array[235] = 32'h00b79023;
    assign array[236] = 32'h05100713;
    assign array[237] = 32'h00e79023;
    assign array[238] = 32'h42100713;
    assign array[239] = 32'h00e79023;
    assign array[240] = 32'h04100713;
    assign array[241] = 32'h00e79023;
    assign array[242] = 32'h00079023;
    assign array[243] = 32'h0037c383;
    assign array[244] = 32'h0037c683;
    assign array[245] = 32'h0037c703;
    assign array[246] = 32'h06e203c2;
    assign array[247] = 32'h00d3e3b3;
    assign array[248] = 32'h0037c683;
    assign array[249] = 32'h0083d393;
    assign array[250] = 32'h67330762;
    assign array[251] = 32'h83210077;
    assign array[252] = 32'h82a306e2;
    assign array[253] = 32'h8f5500c7;
    assign array[254] = 32'h00e28a63;
    assign array[255] = 32'h464157b7;
    assign array[256] = 32'h70000737;
    assign array[257] = 32'h94c78793;
    assign array[258] = 32'ha001c31c;
    assign array[259] = 32'h00435683;
    assign array[260] = 32'h00c78223;
    assign array[261] = 32'h00a78123;
    assign array[262] = 32'h00b79023;
    assign array[263] = 32'h600007b7;
    assign array[264] = 32'h0007d703;
    assign array[265] = 32'hff6d8b09;
    assign array[266] = 32'h00078123;
    assign array[267] = 32'h00078123;
    assign array[268] = 32'h81234711;
    assign array[269] = 32'h071300e7;
    assign array[270] = 32'h90230510;
    assign array[271] = 32'h073700e7;
    assign array[272] = 32'h57836000;
    assign array[273] = 32'h8b890007;
    assign array[274] = 32'h0793ffed;
    assign array[275] = 32'h10234210;
    assign array[276] = 32'h07b700f7;
    assign array[277] = 32'hd7036000;
    assign array[278] = 32'h8b090007;
    assign array[279] = 32'h4709ff6d;
    assign array[280] = 32'h00e782a3;
    assign array[281] = 32'h04100713;
    assign array[282] = 32'h00e79023;
    assign array[283] = 32'h60000737;
    assign array[284] = 32'h00075783;
    assign array[285] = 32'hffed8b89;
    assign array[286] = 32'h00071023;
    assign array[287] = 32'h00374603;
    assign array[288] = 32'h00374783;
    assign array[289] = 32'h02a34589;
    assign array[290] = 32'h07a200b7;
    assign array[291] = 32'h8a638fd1;
    assign array[292] = 32'h57b700f6;
    assign array[293] = 32'h07374641;
    assign array[294] = 32'h87937000;
    assign array[295] = 32'hc31c94c7;
    assign array[296] = 32'h8082a001;
    assign array[297] = 32'h07b7671d;
    assign array[298] = 32'h07136000;
    assign array[299] = 32'h9323b827;
    assign array[300] = 32'h460900e7;
    assign array[301] = 32'h30000337;
    assign array[302] = 32'h00032283;
    assign array[303] = 32'h00c78223;
    assign array[304] = 32'h00c782a3;
    assign array[305] = 32'h06b00513;
    assign array[306] = 32'h00a78123;
    assign array[307] = 32'h00078123;
    assign array[308] = 32'h00078123;
    assign array[309] = 32'h00078123;
    assign array[310] = 32'h11100593;
    assign array[311] = 32'h00b79023;
    assign array[312] = 32'h90234745;
    assign array[313] = 32'h670500e7;
    assign array[314] = 32'h82170713;
    assign array[315] = 32'h00e79023;
    assign array[316] = 32'h08100713;
    assign array[317] = 32'h00e79023;
    assign array[318] = 32'h00079023;
    assign array[319] = 32'h0037c383;
    assign array[320] = 32'h0037c683;
    assign array[321] = 32'h0037c703;
    assign array[322] = 32'h06e203c2;
    assign array[323] = 32'h00d3e3b3;
    assign array[324] = 32'h0037c683;
    assign array[325] = 32'h0083d393;
    assign array[326] = 32'h67330762;
    assign array[327] = 32'h83210077;
    assign array[328] = 32'h82a306e2;
    assign array[329] = 32'h8f5500c7;
    assign array[330] = 32'h00e28a63;
    assign array[331] = 32'h464157b7;
    assign array[332] = 32'h70000737;
    assign array[333] = 32'h94c78793;
    assign array[334] = 32'ha001c31c;
    assign array[335] = 32'h00435683;
    assign array[336] = 32'h00c78223;
    assign array[337] = 32'h00a78123;
    assign array[338] = 32'h00b79023;
    assign array[339] = 32'h600007b7;
    assign array[340] = 32'h0007d703;
    assign array[341] = 32'hff6d8b09;
    assign array[342] = 32'h00078123;
    assign array[343] = 32'h00078123;
    assign array[344] = 32'h81234711;
    assign array[345] = 32'h474500e7;
    assign array[346] = 32'h00e79023;
    assign array[347] = 32'h60000737;
    assign array[348] = 32'h00075783;
    assign array[349] = 32'hffed8b89;
    assign array[350] = 32'h87936785;
    assign array[351] = 32'h10238217;
    assign array[352] = 32'h07b700f7;
    assign array[353] = 32'hd7036000;
    assign array[354] = 32'h8b090007;
    assign array[355] = 32'h4709ff6d;
    assign array[356] = 32'h00e782a3;
    assign array[357] = 32'h08100713;
    assign array[358] = 32'h00e79023;
    assign array[359] = 32'h60000737;
    assign array[360] = 32'h00075783;
    assign array[361] = 32'hffed8b89;
    assign array[362] = 32'h00071023;
    assign array[363] = 32'h00374603;
    assign array[364] = 32'h00374783;
    assign array[365] = 32'h02a34589;
    assign array[366] = 32'h07a200b7;
    assign array[367] = 32'h8a638fd1;
    assign array[368] = 32'h57b700f6;
    assign array[369] = 32'h07374641;
    assign array[370] = 32'h87937000;
    assign array[371] = 32'hc31c94c7;
    assign array[372] = 32'h8082a001;
    assign array[373] = 32'h07b7777d;
    assign array[374] = 32'h07136000;
    assign array[375] = 32'h9323b647;
    assign array[376] = 32'h460900e7;
    assign array[377] = 32'h30000337;
    assign array[378] = 32'h00032283;
    assign array[379] = 32'h00c78223;
    assign array[380] = 32'h00c782a3;
    assign array[381] = 32'h8123552d;
    assign array[382] = 32'h812300a7;
    assign array[383] = 32'h81230007;
    assign array[384] = 32'h81230007;
    assign array[385] = 32'h05930007;
    assign array[386] = 32'h90231110;
    assign array[387] = 32'h071300b7;
    assign array[388] = 32'h90230910;
    assign array[389] = 32'h071300e7;
    assign array[390] = 32'h90236210;
    assign array[391] = 32'h071300e7;
    assign array[392] = 32'h90230810;
    assign array[393] = 32'h902300e7;
    assign array[394] = 32'hc3830007;
    assign array[395] = 32'hc6830037;
    assign array[396] = 32'hc7030037;
    assign array[397] = 32'h03c20037;
    assign array[398] = 32'he3b306e2;
    assign array[399] = 32'hc68300d3;
    assign array[400] = 32'hd3930037;
    assign array[401] = 32'h07620083;
    assign array[402] = 32'h00776733;
    assign array[403] = 32'h06e28321;
    assign array[404] = 32'h00c782a3;
    assign array[405] = 32'h8a638f55;
    assign array[406] = 32'h57b700e2;
    assign array[407] = 32'h07374641;
    assign array[408] = 32'h87937000;
    assign array[409] = 32'hc31c94c7;
    assign array[410] = 32'h5683a001;
    assign array[411] = 32'h82230043;
    assign array[412] = 32'h812300c7;
    assign array[413] = 32'h902300a7;
    assign array[414] = 32'h07b700b7;
    assign array[415] = 32'hd7036000;
    assign array[416] = 32'h8b090007;
    assign array[417] = 32'h8123ff6d;
    assign array[418] = 32'h81230007;
    assign array[419] = 32'h47110007;
    assign array[420] = 32'h00e78123;
    assign array[421] = 32'h09100713;
    assign array[422] = 32'h00e79023;
    assign array[423] = 32'h60000737;
    assign array[424] = 32'h00075783;
    assign array[425] = 32'hffed8b89;
    assign array[426] = 32'h62100793;
    assign array[427] = 32'h00f71023;
    assign array[428] = 32'h600007b7;
    assign array[429] = 32'h0007d703;
    assign array[430] = 32'hff6d8b09;
    assign array[431] = 32'h82a34709;
    assign array[432] = 32'h071300e7;
    assign array[433] = 32'h90230810;
    assign array[434] = 32'h073700e7;
    assign array[435] = 32'h57836000;
    assign array[436] = 32'h8b890007;
    assign array[437] = 32'h1023ffed;
    assign array[438] = 32'h46030007;
    assign array[439] = 32'h47830037;
    assign array[440] = 32'h45890037;
    assign array[441] = 32'h00b702a3;
    assign array[442] = 32'h8fd107a2;
    assign array[443] = 32'h00f68a63;
    assign array[444] = 32'h464157b7;
    assign array[445] = 32'h70000737;
    assign array[446] = 32'h94c78793;
    assign array[447] = 32'ha001c31c;
    assign array[448] = 32'h77718082;
    assign array[449] = 32'h600007b7;
    assign array[450] = 32'hb8570713;
    assign array[451] = 32'h00e79323;
    assign array[452] = 32'h03374609;
    assign array[453] = 32'h22833000;
    assign array[454] = 32'h82230003;
    assign array[455] = 32'h82a300c7;
    assign array[456] = 32'h051300c7;
    assign array[457] = 32'h8123fbb0;
    assign array[458] = 32'h812300a7;
    assign array[459] = 32'h81230007;
    assign array[460] = 32'h81230007;
    assign array[461] = 32'h05930007;
    assign array[462] = 32'h90231510;
    assign array[463] = 32'h071300b7;
    assign array[464] = 32'h90230510;
    assign array[465] = 32'h670500e7;
    assign array[466] = 32'h82170713;
    assign array[467] = 32'h00e79023;
    assign array[468] = 32'h04100713;
    assign array[469] = 32'h00e79023;
    assign array[470] = 32'h00079023;
    assign array[471] = 32'h0037c383;
    assign array[472] = 32'h0037c683;
    assign array[473] = 32'h0037c703;
    assign array[474] = 32'h06e203c2;
    assign array[475] = 32'h00d3e3b3;
    assign array[476] = 32'h0037c683;
    assign array[477] = 32'h0083d393;
    assign array[478] = 32'h67330762;
    assign array[479] = 32'h83210077;
    assign array[480] = 32'h82a306e2;
    assign array[481] = 32'h8f5500c7;
    assign array[482] = 32'h00e28a63;
    assign array[483] = 32'h464157b7;
    assign array[484] = 32'h70000737;
    assign array[485] = 32'h94c78793;
    assign array[486] = 32'ha001c31c;
    assign array[487] = 32'h00435683;
    assign array[488] = 32'h00c78223;
    assign array[489] = 32'h00a78123;
    assign array[490] = 32'h00b79023;
    assign array[491] = 32'h600007b7;
    assign array[492] = 32'h0007d703;
    assign array[493] = 32'hff6d8b09;
    assign array[494] = 32'h00078123;
    assign array[495] = 32'h00078123;
    assign array[496] = 32'h81234711;
    assign array[497] = 32'h071300e7;
    assign array[498] = 32'h90230510;
    assign array[499] = 32'h073700e7;
    assign array[500] = 32'h57836000;
    assign array[501] = 32'h8b890007;
    assign array[502] = 32'h6785ffed;
    assign array[503] = 32'h82178793;
    assign array[504] = 32'h00f71023;
    assign array[505] = 32'h600007b7;
    assign array[506] = 32'h0007d703;
    assign array[507] = 32'hff6d8b09;
    assign array[508] = 32'h82a34709;
    assign array[509] = 32'h071300e7;
    assign array[510] = 32'h90230410;
    assign array[511] = 32'h073700e7;
    assign array[512] = 32'h57836000;
    assign array[513] = 32'h8b890007;
    assign array[514] = 32'h1023ffed;
    assign array[515] = 32'h46030007;
    assign array[516] = 32'h47830037;
    assign array[517] = 32'h45890037;
    assign array[518] = 32'h00b702a3;
    assign array[519] = 32'h8fd107a2;
    assign array[520] = 32'h00f68a63;
    assign array[521] = 32'h464157b7;
    assign array[522] = 32'h70000737;
    assign array[523] = 32'h94c78793;
    assign array[524] = 32'ha001c31c;
    assign array[525] = 32'h777d8082;
    assign array[526] = 32'h600007b7;
    assign array[527] = 32'hba670713;
    assign array[528] = 32'h00e79323;
    assign array[529] = 32'h03374609;
    assign array[530] = 32'h22833000;
    assign array[531] = 32'h82230003;
    assign array[532] = 32'h82a300c7;
    assign array[533] = 32'h552d00c7;
    assign array[534] = 32'h00a78123;
    assign array[535] = 32'h00078123;
    assign array[536] = 32'h00078123;
    assign array[537] = 32'h00078123;
    assign array[538] = 32'h19100593;
    assign array[539] = 32'h00b79023;
    assign array[540] = 32'h09100713;
    assign array[541] = 32'h00e79023;
    assign array[542] = 32'h07136705;
    assign array[543] = 32'h9023a217;
    assign array[544] = 32'h071300e7;
    assign array[545] = 32'h90230810;
    assign array[546] = 32'h902300e7;
    assign array[547] = 32'hc3830007;
    assign array[548] = 32'hc6830037;
    assign array[549] = 32'hc7030037;
    assign array[550] = 32'h03c20037;
    assign array[551] = 32'he3b306e2;
    assign array[552] = 32'hc68300d3;
    assign array[553] = 32'hd3930037;
    assign array[554] = 32'h07620083;
    assign array[555] = 32'h00776733;
    assign array[556] = 32'h06e28321;
    assign array[557] = 32'h00c782a3;
    assign array[558] = 32'h8a638f55;
    assign array[559] = 32'h57b700e2;
    assign array[560] = 32'h07374641;
    assign array[561] = 32'h87937000;
    assign array[562] = 32'hc31c94c7;
    assign array[563] = 32'h5683a001;
    assign array[564] = 32'h82230043;
    assign array[565] = 32'h812300c7;
    assign array[566] = 32'h902300a7;
    assign array[567] = 32'h07b700b7;
    assign array[568] = 32'hd7036000;
    assign array[569] = 32'h8b090007;
    assign array[570] = 32'h8123ff6d;
    assign array[571] = 32'h81230007;
    assign array[572] = 32'h47110007;
    assign array[573] = 32'h00e78123;
    assign array[574] = 32'h09100713;
    assign array[575] = 32'h00e79023;
    assign array[576] = 32'h60000737;
    assign array[577] = 32'h00075783;
    assign array[578] = 32'hffed8b89;
    assign array[579] = 32'h87936785;
    assign array[580] = 32'h1023a217;
    assign array[581] = 32'h07b700f7;
    assign array[582] = 32'hd7036000;
    assign array[583] = 32'h8b090007;
    assign array[584] = 32'h4709ff6d;
    assign array[585] = 32'h00e782a3;
    assign array[586] = 32'h08100713;
    assign array[587] = 32'h00e79023;
    assign array[588] = 32'h60000737;
    assign array[589] = 32'h00075783;
    assign array[590] = 32'hffed8b89;
    assign array[591] = 32'h00071023;
    assign array[592] = 32'h00374603;
    assign array[593] = 32'h00374783;
    assign array[594] = 32'h02a34589;
    assign array[595] = 32'h07a200b7;
    assign array[596] = 32'h8a638fd1;
    assign array[597] = 32'h57b700f6;
    assign array[598] = 32'h07374641;
    assign array[599] = 32'h87937000;
    assign array[600] = 32'hc31c94c7;
    assign array[601] = 32'h8082a001;
    assign array[602] = 32'h57b71151;
    assign array[603] = 32'hc4065153;
    assign array[604] = 32'h04978793;
    assign array[605] = 32'h0437c222;
    assign array[606] = 32'hc01c7000;
    assign array[607] = 32'he98ff0ef;
    assign array[608] = 32'hf9cff0ef;
    assign array[609] = 32'h32fd30c1;
    assign array[610] = 32'h31a93e31;
    assign array[611] = 32'h443257b7;
    assign array[612] = 32'h04978793;
    assign array[613] = 32'h33b5c01c;
    assign array[614] = 32'h513457b7;
    assign array[615] = 32'h04978793;
    assign array[616] = 32'h3d51c01c;
    assign array[617] = 32'h504157b7;
    assign array[618] = 32'h35378793;
    assign array[619] = 32'ha001c01c;
    assign array[620] = 32'h00000014;
    assign array[621] = 32'h00000000;
    assign array[622] = 32'h00527a01;
    assign array[623] = 32'h01017c01;
    assign array[624] = 32'h07020d1b;
    assign array[625] = 32'h00000001;
    assign array[626] = 32'h00000010;
    assign array[627] = 32'h0000001c;
    assign array[628] = 32'hfffff630;
    assign array[629] = 32'h00000014;
    assign array[630] = 32'h00000000;
