    assign array[0] = 32'h10001197;
    assign array[1] = 32'h80018193;
    assign array[2] = 32'h10000117;
    assign array[3] = 32'h1f810113;
    assign array[4] = 32'h1171203d;
    assign array[5] = 32'h0040c022;
    assign array[6] = 32'h700007b7;
    assign array[7] = 32'h50415737;
    assign array[8] = 32'h35370713;
    assign array[9] = 32'ha001c398;
    assign array[10] = 32'hc0221171;
    assign array[11] = 32'h07b70040;
    assign array[12] = 32'h57377000;
    assign array[13] = 32'h07134641;
    assign array[14] = 32'hc39894c7;
    assign array[15] = 32'h1121a001;
    assign array[16] = 32'hc822ca06;
    assign array[17] = 32'h07b70820;
    assign array[18] = 32'h07136000;
    assign array[19] = 32'h93233000;
    assign array[20] = 32'h07b700e7;
    assign array[21] = 32'h439c3000;
    assign array[22] = 32'hfef42823;
    assign array[23] = 32'h600007b7;
    assign array[24] = 32'h82234709;
    assign array[25] = 32'h07b700e7;
    assign array[26] = 32'h470d6000;
    assign array[27] = 32'h00e78123;
    assign array[28] = 32'h600007b7;
    assign array[29] = 32'h10500713;
    assign array[30] = 32'h00e79023;
    assign array[31] = 32'h600007b7;
    assign array[32] = 32'h00078123;
    assign array[33] = 32'h600007b7;
    assign array[34] = 32'h00078123;
    assign array[35] = 32'h600007b7;
    assign array[36] = 32'h00078123;
    assign array[37] = 32'h600007b7;
    assign array[38] = 32'h90234715;
    assign array[39] = 32'h07b700e7;
    assign array[40] = 32'h47096000;
    assign array[41] = 32'h00e782a3;
    assign array[42] = 32'h600007b7;
    assign array[43] = 32'h90234705;
    assign array[44] = 32'h07b700e7;
    assign array[45] = 32'h90236000;
    assign array[46] = 32'h26230007;
    assign array[47] = 32'h07b7fe04;
    assign array[48] = 32'hc7836000;
    assign array[49] = 32'hf7930037;
    assign array[50] = 32'h07e20ff7;
    assign array[51] = 32'h2783873e;
    assign array[52] = 32'h83a1fec4;
    assign array[53] = 32'h26238fd9;
    assign array[54] = 32'h07b7fef4;
    assign array[55] = 32'hc7836000;
    assign array[56] = 32'hf7930037;
    assign array[57] = 32'h07e20ff7;
    assign array[58] = 32'h2783873e;
    assign array[59] = 32'h83a1fec4;
    assign array[60] = 32'h26238fd9;
    assign array[61] = 32'h07b7fef4;
    assign array[62] = 32'hc7836000;
    assign array[63] = 32'hf7930037;
    assign array[64] = 32'h07e20ff7;
    assign array[65] = 32'h2783873e;
    assign array[66] = 32'h83a1fec4;
    assign array[67] = 32'h26238fd9;
    assign array[68] = 32'h07b7fef4;
    assign array[69] = 32'hc7836000;
    assign array[70] = 32'hf7930037;
    assign array[71] = 32'h07e20ff7;
    assign array[72] = 32'h2783873e;
    assign array[73] = 32'h83a1fec4;
    assign array[74] = 32'h26238fd9;
    assign array[75] = 32'h07b7fef4;
    assign array[76] = 32'h47096000;
    assign array[77] = 32'h00e782a3;
    assign array[78] = 32'hff042703;
    assign array[79] = 32'hfec42783;
    assign array[80] = 32'h00f70363;
    assign array[81] = 32'h07b735d5;
    assign array[82] = 32'h07913000;
    assign array[83] = 32'h0007d783;
    assign array[84] = 32'hfef41523;
    assign array[85] = 32'h600007b7;
    assign array[86] = 32'h82234709;
    assign array[87] = 32'h07b700e7;
    assign array[88] = 32'h470d6000;
    assign array[89] = 32'h00e78123;
    assign array[90] = 32'h600007b7;
    assign array[91] = 32'h10500713;
    assign array[92] = 32'h00e79023;
    assign array[93] = 32'h600007b7;
    assign array[94] = 32'h00078123;
    assign array[95] = 32'h600007b7;
    assign array[96] = 32'h00078123;
    assign array[97] = 32'h600007b7;
    assign array[98] = 32'h81234711;
    assign array[99] = 32'h07b700e7;
    assign array[100] = 32'h47156000;
    assign array[101] = 32'h00e79023;
    assign array[102] = 32'h600007b7;
    assign array[103] = 32'h82a34709;
    assign array[104] = 32'h07b700e7;
    assign array[105] = 32'h47056000;
    assign array[106] = 32'h00e79023;
    assign array[107] = 32'h600007b7;
    assign array[108] = 32'h00079023;
    assign array[109] = 32'hfe041423;
    assign array[110] = 32'h600007b7;
    assign array[111] = 32'h0037c783;
    assign array[112] = 32'h0ff7f793;
    assign array[113] = 32'h971307a2;
    assign array[114] = 32'h87410107;
    assign array[115] = 32'hfe845783;
    assign array[116] = 32'h07c283a1;
    assign array[117] = 32'h07c283c1;
    assign array[118] = 32'h8fd987c1;
    assign array[119] = 32'h87c107c2;
    assign array[120] = 32'hfef41423;
    assign array[121] = 32'h600007b7;
    assign array[122] = 32'h0037c783;
    assign array[123] = 32'h0ff7f793;
    assign array[124] = 32'h971307a2;
    assign array[125] = 32'h87410107;
    assign array[126] = 32'hfe845783;
    assign array[127] = 32'h07c283a1;
    assign array[128] = 32'h07c283c1;
    assign array[129] = 32'h8fd987c1;
    assign array[130] = 32'h87c107c2;
    assign array[131] = 32'hfef41423;
    assign array[132] = 32'h600007b7;
    assign array[133] = 32'h82a34709;
    assign array[134] = 32'h07b700e7;
    assign array[135] = 32'h57037000;
    assign array[136] = 32'hc398fea4;
    assign array[137] = 32'h700007b7;
    assign array[138] = 32'hfe845703;
    assign array[139] = 32'h5703c398;
    assign array[140] = 32'h5783fea4;
    assign array[141] = 32'h0363fe84;
    assign array[142] = 32'h33fd00f7;
    assign array[143] = 32'h47813bd9;
    assign array[144] = 32'h40d2853e;
    assign array[145] = 32'h01614442;
    assign array[146] = 32'h00008082;
    assign array[147] = 32'h00000014;
    assign array[148] = 32'h00000000;
    assign array[149] = 32'h00527a01;
    assign array[150] = 32'h01017c01;
    assign array[151] = 32'h07020d1b;
    assign array[152] = 32'h00000001;
    assign array[153] = 32'h00000010;
    assign array[154] = 32'h0000001c;
    assign array[155] = 32'hfffffd94;
    assign array[156] = 32'h00000012;
    assign array[157] = 32'h00000000;
