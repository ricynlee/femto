    assign array[0] = 32'h10001197;
    assign array[1] = 32'h80018193;
    assign array[2] = 32'h10000117;
    assign array[3] = 32'h1f810113;
    assign array[4] = 32'h11712015;
    assign array[5] = 32'h0040c022;
    assign array[6] = 32'hf00007b7;
    assign array[7] = 32'h00078023;
    assign array[8] = 32'h1171a001;
    assign array[9] = 32'h0040c022;
    assign array[10] = 32'hf00007b7;
    assign array[11] = 32'h80234705;
    assign array[12] = 32'ha00100e7;
    assign array[13] = 32'hc4061151;
    assign array[14] = 32'h0060c222;
    assign array[15] = 32'h200007b7;
    assign array[16] = 32'h0793873e;
    assign array[17] = 32'h002305a0;
    assign array[18] = 32'h07b700f7;
    assign array[19] = 32'hc7032000;
    assign array[20] = 32'h07930007;
    assign array[21] = 32'h036305a0;
    assign array[22] = 32'h37e100f7;
    assign array[23] = 32'h200007b7;
    assign array[24] = 32'h6799873e;
    assign array[25] = 32'ha3c78793;
    assign array[26] = 32'h00f71023;
    assign array[27] = 32'h200007b7;
    assign array[28] = 32'h0007d703;
    assign array[29] = 32'h87936799;
    assign array[30] = 32'h0363a3c7;
    assign array[31] = 32'h375500f7;
    assign array[32] = 32'h200007b7;
    assign array[33] = 32'h77b7873e;
    assign array[34] = 32'h87935a3c;
    assign array[35] = 32'hc31c92d7;
    assign array[36] = 32'h200007b7;
    assign array[37] = 32'h77b74398;
    assign array[38] = 32'h87935a3c;
    assign array[39] = 32'h036392d7;
    assign array[40] = 32'h374100f7;
    assign array[41] = 32'h478137bd;
    assign array[42] = 32'h40a2853e;
    assign array[43] = 32'h01314412;
    assign array[44] = 32'h00008082;
    assign array[45] = 32'h00000014;
    assign array[46] = 32'h00000000;
    assign array[47] = 32'h00527a01;
    assign array[48] = 32'h01017c01;
    assign array[49] = 32'h07020d1b;
    assign array[50] = 32'h00000001;
    assign array[51] = 32'h00000010;
    assign array[52] = 32'h0000001c;
    assign array[53] = 32'hffffff2c;
    assign array[54] = 32'h00000012;
    assign array[55] = 32'h00000000;
    assign array[56] = 32'h20000000;
