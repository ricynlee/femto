    assign array[0] = 8'h97;
    assign array[1] = 8'h11;
    assign array[2] = 8'hd4;
    assign array[3] = 8'hef;
    assign array[4] = 8'h93;
    assign array[5] = 8'h81;
    assign array[6] = 8'h01;
    assign array[7] = 8'h80;
    assign array[8] = 8'h17;
    assign array[9] = 8'h01;
    assign array[10] = 8'hd4;
    assign array[11] = 8'hef;
    assign array[12] = 8'h13;
    assign array[13] = 8'h01;
    assign array[14] = 8'h81;
    assign array[15] = 8'h1f;
    assign array[16] = 8'hef;
    assign array[17] = 8'h00;
    assign array[18] = 8'h40;
    assign array[19] = 8'h00;
    assign array[20] = 8'h13;
    assign array[21] = 8'h01;
    assign array[22] = 8'h81;
    assign array[23] = 8'hff;
    assign array[24] = 8'h23;
    assign array[25] = 8'h22;
    assign array[26] = 8'h81;
    assign array[27] = 8'h00;
    assign array[28] = 8'h13;
    assign array[29] = 8'h04;
    assign array[30] = 8'h81;
    assign array[31] = 8'h00;
    assign array[32] = 8'hb7;
    assign array[33] = 8'h07;
    assign array[34] = 8'h00;
    assign array[35] = 8'h40;
    assign array[36] = 8'h13;
    assign array[37] = 8'h07;
    assign array[38] = 8'h80;
    assign array[39] = 8'h00;
    assign array[40] = 8'h23;
    assign array[41] = 8'ha2;
    assign array[42] = 8'he7;
    assign array[43] = 8'h00;
    assign array[44] = 8'hb7;
    assign array[45] = 8'h07;
    assign array[46] = 8'h00;
    assign array[47] = 8'h40;
    assign array[48] = 8'h13;
    assign array[49] = 8'h07;
    assign array[50] = 8'h80;
    assign array[51] = 8'h00;
    assign array[52] = 8'h23;
    assign array[53] = 8'ha0;
    assign array[54] = 8'he7;
    assign array[55] = 8'h00;
    assign array[56] = 8'h23;
    assign array[57] = 8'h2c;
    assign array[58] = 8'h04;
    assign array[59] = 8'hfe;
    assign array[60] = 8'h6f;
    assign array[61] = 8'h00;
    assign array[62] = 8'h00;
    assign array[63] = 8'h01;
    assign array[64] = 8'h83;
    assign array[65] = 8'h27;
    assign array[66] = 8'h84;
    assign array[67] = 8'hff;
    assign array[68] = 8'h93;
    assign array[69] = 8'h87;
    assign array[70] = 8'h17;
    assign array[71] = 8'h00;
    assign array[72] = 8'h23;
    assign array[73] = 8'h2c;
    assign array[74] = 8'hf4;
    assign array[75] = 8'hfe;
    assign array[76] = 8'h03;
    assign array[77] = 8'h27;
    assign array[78] = 8'h84;
    assign array[79] = 8'hff;
    assign array[80] = 8'hb7;
    assign array[81] = 8'h17;
    assign array[82] = 8'h00;
    assign array[83] = 8'h00;
    assign array[84] = 8'h93;
    assign array[85] = 8'h87;
    assign array[86] = 8'h77;
    assign array[87] = 8'h38;
    assign array[88] = 8'he3;
    assign array[89] = 8'hd4;
    assign array[90] = 8'he7;
    assign array[91] = 8'hfe;
    assign array[92] = 8'hb7;
    assign array[93] = 8'h07;
    assign array[94] = 8'h00;
    assign array[95] = 8'h40;
    assign array[96] = 8'h03;
    assign array[97] = 8'ha7;
    assign array[98] = 8'h07;
    assign array[99] = 8'h00;
    assign array[100] = 8'hb7;
    assign array[101] = 8'h07;
    assign array[102] = 8'h00;
    assign array[103] = 8'h40;
    assign array[104] = 8'h13;
    assign array[105] = 8'h47;
    assign array[106] = 8'h87;
    assign array[107] = 8'h00;
    assign array[108] = 8'h23;
    assign array[109] = 8'ha0;
    assign array[110] = 8'he7;
    assign array[111] = 8'h00;
    assign array[112] = 8'h6f;
    assign array[113] = 8'hf0;
    assign array[114] = 8'h9f;
    assign array[115] = 8'hfc;
    assign array[116] = 8'h14;
    assign array[117] = 8'h00;
    assign array[118] = 8'h00;
    assign array[119] = 8'h00;
    assign array[120] = 8'h00;
    assign array[121] = 8'h00;
    assign array[122] = 8'h00;
    assign array[123] = 8'h00;
    assign array[124] = 8'h01;
    assign array[125] = 8'h7a;
    assign array[126] = 8'h52;
    assign array[127] = 8'h00;
    assign array[128] = 8'h01;
    assign array[129] = 8'h7c;
    assign array[130] = 8'h01;
    assign array[131] = 8'h01;
    assign array[132] = 8'h1b;
    assign array[133] = 8'h0d;
    assign array[134] = 8'h02;
    assign array[135] = 8'h07;
    assign array[136] = 8'h01;
    assign array[137] = 8'h00;
    assign array[138] = 8'h00;
    assign array[139] = 8'h00;
    assign array[140] = 8'h10;
    assign array[141] = 8'h00;
    assign array[142] = 8'h00;
    assign array[143] = 8'h00;
    assign array[144] = 8'h1c;
    assign array[145] = 8'h00;
    assign array[146] = 8'h00;
    assign array[147] = 8'h00;
    assign array[148] = 8'h6c;
    assign array[149] = 8'hff;
    assign array[150] = 8'hff;
    assign array[151] = 8'hff;
    assign array[152] = 8'h14;
    assign array[153] = 8'h00;
    assign array[154] = 8'h00;
    assign array[155] = 8'h00;
    assign array[156] = 8'h00;
    assign array[157] = 8'h00;
    assign array[158] = 8'h00;
    assign array[159] = 8'h00;
    assign array[160] = 8'h00;
    assign array[161] = 8'h00;
    assign array[162] = 8'h00;
    assign array[163] = 8'h40;
    assign array[164] = 8'h00;
    assign array[165] = 8'h00;
    assign array[166] = 8'h00;
    assign array[167] = 8'h50;
