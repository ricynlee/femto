module ioring();

endmodule
