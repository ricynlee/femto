    assign array[0] = 32'h10001197;
    assign array[1] = 32'h80018193;
    assign array[2] = 32'h10000117;
    assign array[3] = 32'h1f810113;
    assign array[4] = 32'h20152019;
    assign array[5] = 32'h06b72889;
    assign array[6] = 32'h07131000;
    assign array[7] = 32'h47810000;
    assign array[8] = 32'h00068693;
    assign array[9] = 32'h00e7e363;
    assign array[10] = 32'h86338082;
    assign array[11] = 32'h002300d7;
    assign array[12] = 32'h07850006;
    assign array[13] = 32'h0637bfc5;
    assign array[14] = 32'h07131000;
    assign array[15] = 32'h47810000;
    assign array[16] = 32'h41c00693;
    assign array[17] = 32'h00060613;
    assign array[18] = 32'h00e7e363;
    assign array[19] = 32'h85b38082;
    assign array[20] = 32'hc58300d7;
    assign array[21] = 32'h85330005;
    assign array[22] = 32'h078500c7;
    assign array[23] = 32'h0ff5f593;
    assign array[24] = 32'h00b50023;
    assign array[25] = 32'h1151b7d5;
    assign array[26] = 32'hc406c222;
    assign array[27] = 32'h20994401;
    assign array[28] = 32'hdd7d2819;
    assign array[29] = 32'hfd7d2809;
    assign array[30] = 32'h46018522;
    assign array[31] = 32'h20314581;
    assign array[32] = 32'h00144413;
    assign array[33] = 32'h4501b7f5;
    assign array[34] = 32'h1141a07d;
    assign array[35] = 32'h842ec422;
    assign array[36] = 32'h00154593;
    assign array[37] = 32'hc6064505;
    assign array[38] = 32'h206dc032;
    assign array[39] = 32'h00144593;
    assign array[40] = 32'h204d4509;
    assign array[41] = 32'h44224602;
    assign array[42] = 32'h459340b2;
    assign array[43] = 32'h450d0016;
    assign array[44] = 32'ha8490141;
    assign array[45] = 32'h46011151;
    assign array[46] = 32'h45014581;
    assign array[47] = 32'h37f1c406;
    assign array[48] = 32'h45014581;
    assign array[49] = 32'h45852881;
    assign array[50] = 32'h20a94505;
    assign array[51] = 32'h45094585;
    assign array[52] = 32'h40a22091;
    assign array[53] = 32'h450d4585;
    assign array[54] = 32'ha82d0131;
    assign array[55] = 32'h02054363;
    assign array[56] = 32'hd3634799;
    assign array[57] = 32'h451900a7;
    assign array[58] = 32'h76130612;
    assign array[59] = 32'h05a20ff6;
    assign array[60] = 32'h8e498e4d;
    assign array[61] = 32'h82410642;
    assign array[62] = 32'h600007b7;
    assign array[63] = 32'h00c79323;
    assign array[64] = 32'h45018082;
    assign array[65] = 32'h07b7b7d5;
    assign array[66] = 32'h43dc4000;
    assign array[67] = 32'h00a7d533;
    assign array[68] = 32'h80828905;
    assign array[69] = 32'h400007b7;
    assign array[70] = 32'h470543dc;
    assign array[71] = 32'h00a71533;
    assign array[72] = 32'h00e59763;
    assign array[73] = 32'h07378fc9;
    assign array[74] = 32'hc35c4000;
    assign array[75] = 32'h45138082;
    assign array[76] = 32'h8fe9fff5;
    assign array[77] = 32'h07b7bfcd;
    assign array[78] = 32'h439c4000;
    assign array[79] = 32'h00a7d533;
    assign array[80] = 32'h80828905;
    assign array[81] = 32'h95334785;
    assign array[82] = 32'hc59900a7;
    assign array[83] = 32'h40000737;
    assign array[84] = 32'h8d5d431c;
    assign array[85] = 32'h8082c308;
    assign array[86] = 32'h400007b7;
    assign array[87] = 32'h45134398;
    assign array[88] = 32'h8d79fff5;
    assign array[89] = 32'h8082c388;
    assign array[90] = 32'hc2221151;
    assign array[91] = 32'h842ac406;
    assign array[92] = 32'h459337d9;
    assign array[93] = 32'h85220015;
    assign array[94] = 32'h40a24412;
    assign array[95] = 32'h0ff5f593;
    assign array[96] = 32'hb7c90131;
    assign array[97] = 32'h500007b7;
    assign array[98] = 32'h0037c503;
    assign array[99] = 32'h80828905;
    assign array[100] = 32'h500007b7;
    assign array[101] = 32'h0027c503;
    assign array[102] = 32'h80828905;
    assign array[103] = 32'h500007b7;
    assign array[104] = 32'h81a34709;
    assign array[105] = 32'h808200e7;
    assign array[106] = 32'h4501e901;
    assign array[107] = 32'h45018082;
    assign array[108] = 32'h441240a2;
    assign array[109] = 32'h80820131;
    assign array[110] = 32'hc2221151;
    assign array[111] = 32'h842ac406;
    assign array[112] = 32'hd57537d1;
    assign array[113] = 32'h500007b7;
    assign array[114] = 32'h0017c783;
    assign array[115] = 32'h00f40023;
    assign array[116] = 32'h1151b7c5;
    assign array[117] = 32'hc406c222;
    assign array[118] = 32'h3f5d842a;
    assign array[119] = 32'h07b7c509;
    assign array[120] = 32'h80235000;
    assign array[121] = 32'h40a20087;
    assign array[122] = 32'h01314412;
    assign array[123] = 32'h11518082;
    assign array[124] = 32'hc026c222;
    assign array[125] = 32'h842ac406;
    assign array[126] = 32'h00b504b3;
    assign array[127] = 32'h00941763;
    assign array[128] = 32'h441240a2;
    assign array[129] = 32'h01314482;
    assign array[130] = 32'h85228082;
    assign array[131] = 32'hdd753f71;
    assign array[132] = 32'hb7ed0405;
    assign array[133] = 32'hc2221151;
    assign array[134] = 32'hc406c026;
    assign array[135] = 32'h04b3842a;
    assign array[136] = 32'h176300b5;
    assign array[137] = 32'h40a20094;
    assign array[138] = 32'h44824412;
    assign array[139] = 32'h80820131;
    assign array[140] = 32'h00044503;
    assign array[141] = 32'hdd6d3f79;
    assign array[142] = 32'hb7e50405;
    assign array[143] = 32'h600007b7;
    assign array[144] = 32'h0057c503;
    assign array[145] = 32'h3533897d;
    assign array[146] = 32'h808200a0;
    assign array[147] = 32'h600007b7;
    assign array[148] = 32'h0047c503;
    assign array[149] = 32'h3533897d;
    assign array[150] = 32'h808200a0;
    assign array[151] = 32'h07b7c519;
    assign array[152] = 32'h07136000;
    assign array[153] = 32'h82a3f800;
    assign array[154] = 32'hc59900e7;
    assign array[155] = 32'h600007b7;
    assign array[156] = 32'hf8000713;
    assign array[157] = 32'h00e78223;
    assign array[158] = 32'he9018082;
    assign array[159] = 32'h80824501;
    assign array[160] = 32'h40a24501;
    assign array[161] = 32'h01314412;
    assign array[162] = 32'h11518082;
    assign array[163] = 32'hc406c222;
    assign array[164] = 32'h376d842a;
    assign array[165] = 32'h07b7d575;
    assign array[166] = 32'hc7836000;
    assign array[167] = 32'h00230037;
    assign array[168] = 32'hb7c500f4;
    assign array[169] = 32'hc2221151;
    assign array[170] = 32'h842ac406;
    assign array[171] = 32'hc5093745;
    assign array[172] = 32'h600007b7;
    assign array[173] = 32'h00878123;
    assign array[174] = 32'h441240a2;
    assign array[175] = 32'h80820131;
    assign array[176] = 32'h600007b7;
    assign array[177] = 32'h0007d503;
    assign array[178] = 32'h89058105;
    assign array[179] = 32'h67858082;
    assign array[180] = 32'hf0078793;
    assign array[181] = 32'h0522059a;
    assign array[182] = 32'hf5938d7d;
    assign array[183] = 32'h8dc90ff5;
    assign array[184] = 32'h0115e593;
    assign array[185] = 32'h600007b7;
    assign array[186] = 32'h00b79023;
    assign array[187] = 32'h67858082;
    assign array[188] = 32'hf0078793;
    assign array[189] = 32'h0522059a;
    assign array[190] = 32'hf5938d7d;
    assign array[191] = 32'h8dc90ff5;
    assign array[192] = 32'h0015e593;
    assign array[193] = 32'h600007b7;
    assign array[194] = 32'h00b79023;
    assign array[195] = 32'h67858082;
    assign array[196] = 32'hf0078793;
    assign array[197] = 32'h0522059a;
    assign array[198] = 32'hf5938d7d;
    assign array[199] = 32'h8dc90ff5;
    assign array[200] = 32'h0315e593;
    assign array[201] = 32'h600007b7;
    assign array[202] = 32'h00b79023;
    assign array[203] = 32'h07b78082;
    assign array[204] = 32'h90236000;
    assign array[205] = 32'h80820007;
    assign array[206] = 32'h06b74781;
    assign array[207] = 32'he3636000;
    assign array[208] = 32'h808200b7;
    assign array[209] = 32'h0056c703;
    assign array[210] = 32'h8b7d862e;
    assign array[211] = 32'h7363973e;
    assign array[212] = 32'h863a00b7;
    assign array[213] = 32'hfec7f5e3;
    assign array[214] = 32'h0036c303;
    assign array[215] = 32'h00f50733;
    assign array[216] = 32'h00230785;
    assign array[217] = 32'hb7fd0067;
    assign array[218] = 32'h06b74781;
    assign array[219] = 32'he3636000;
    assign array[220] = 32'h808200b7;
    assign array[221] = 32'h0046c703;
    assign array[222] = 32'h8b7d862e;
    assign array[223] = 32'h7363973e;
    assign array[224] = 32'h863a00b7;
    assign array[225] = 32'hfec7f5e3;
    assign array[226] = 32'h00f50733;
    assign array[227] = 32'h00074703;
    assign array[228] = 32'h81230785;
    assign array[229] = 32'hb7fd00e6;
    assign array[230] = 32'h700007b7;
    assign array[231] = 32'h8082c388;
    assign array[232] = 32'h700007b7;
    assign array[233] = 32'h80824388;
    assign array[234] = 32'hf00007b7;
    assign array[235] = 32'h00078023;
    assign array[236] = 32'h07b78082;
    assign array[237] = 32'h4705f000;
    assign array[238] = 32'h00e78023;
    assign array[239] = 32'h07b78082;
    assign array[240] = 32'h471df000;
    assign array[241] = 32'h00e78023;
    assign array[242] = 32'h07b78082;
    assign array[243] = 32'h4719f000;
    assign array[244] = 32'h00e78023;
    assign array[245] = 32'h07b78082;
    assign array[246] = 32'h4721f000;
    assign array[247] = 32'h00e78023;
    assign array[248] = 32'h07b78082;
    assign array[249] = 32'h4725f000;
    assign array[250] = 32'h00e78023;
    assign array[251] = 32'h00008082;
    assign array[252] = 32'h00000014;
    assign array[253] = 32'h00000000;
    assign array[254] = 32'h00527a01;
    assign array[255] = 32'h01017c01;
    assign array[256] = 32'h07020d1b;
    assign array[257] = 32'h00000001;
    assign array[258] = 32'h00000010;
    assign array[259] = 32'h0000001c;
    assign array[260] = 32'hfffffbf0;
    assign array[261] = 32'h00000016;
    assign array[262] = 32'h00000000;
