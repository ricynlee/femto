    assign array[0] = 32'h10001197;
    assign array[1] = 32'h80018193;
    assign array[2] = 32'h10000117;
    assign array[3] = 32'h1f810113;
    assign array[4] = 32'h1171203d;
    assign array[5] = 32'h0040c022;
    assign array[6] = 32'h700007b7;
    assign array[7] = 32'h50415737;
    assign array[8] = 32'h35370713;
    assign array[9] = 32'ha001c398;
    assign array[10] = 32'hc0221171;
    assign array[11] = 32'h07b70040;
    assign array[12] = 32'h57377000;
    assign array[13] = 32'h07134641;
    assign array[14] = 32'hc39894c7;
    assign array[15] = 32'h1131a001;
    assign array[16] = 32'hc622c806;
    assign array[17] = 32'h07b70840;
    assign array[18] = 32'h07137000;
    assign array[19] = 32'hc3981000;
    assign array[20] = 32'h700007b7;
    assign array[21] = 32'h2823439c;
    assign array[22] = 32'h0793fef4;
    assign array[23] = 32'h27031000;
    assign array[24] = 32'h6363ff04;
    assign array[25] = 32'h37c900f7;
    assign array[26] = 32'h700007b7;
    assign array[27] = 32'h2623439c;
    assign array[28] = 32'h2703fef4;
    assign array[29] = 32'h2783fec4;
    assign array[30] = 32'h6363ff04;
    assign array[31] = 32'h376d00f7;
    assign array[32] = 32'h07b70001;
    assign array[33] = 32'h439c7000;
    assign array[34] = 32'h3761ffed;
    assign array[35] = 32'h853e4781;
    assign array[36] = 32'h443240c2;
    assign array[37] = 32'h80820151;
    assign array[38] = 32'h00000014;
    assign array[39] = 32'h00000000;
    assign array[40] = 32'h00527a01;
    assign array[41] = 32'h01017c01;
    assign array[42] = 32'h07020d1b;
    assign array[43] = 32'h00000001;
    assign array[44] = 32'h00000010;
    assign array[45] = 32'h0000001c;
    assign array[46] = 32'hffffff48;
    assign array[47] = 32'h00000012;
    assign array[48] = 32'h00000000;
    assign array[49] = 32'h00000100;
