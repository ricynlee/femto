`define HEX_PATH "D:/Projects/femto/rtl/sim/" 
