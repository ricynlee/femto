    assign array[0] = 32'h10001197;
    assign array[1] = 32'h80018193;
    assign array[2] = 32'h10000117;
    assign array[3] = 32'h1f810113;
    assign array[4] = 32'h20152019;
    assign array[5] = 32'h06b728c1;
    assign array[6] = 32'h07131000;
    assign array[7] = 32'h47810000;
    assign array[8] = 32'h00068693;
    assign array[9] = 32'h00e7e363;
    assign array[10] = 32'h86338082;
    assign array[11] = 32'h002300d7;
    assign array[12] = 32'h07850006;
    assign array[13] = 32'h6685bfc5;
    assign array[14] = 32'h10000637;
    assign array[15] = 32'h00000713;
    assign array[16] = 32'h86934781;
    assign array[17] = 32'h06138606;
    assign array[18] = 32'he3630006;
    assign array[19] = 32'h808200e7;
    assign array[20] = 32'h00d785b3;
    assign array[21] = 32'h0005c583;
    assign array[22] = 32'h00c78533;
    assign array[23] = 32'hf5930785;
    assign array[24] = 32'h00230ff5;
    assign array[25] = 32'hb7d500b5;
    assign array[26] = 32'hc2221151;
    assign array[27] = 32'h440dc406;
    assign array[28] = 32'h45854601;
    assign array[29] = 32'h00ef4501;
    assign array[30] = 32'h053776c0;
    assign array[31] = 32'h2ba50004;
    assign array[32] = 32'h45814601;
    assign array[33] = 32'h00ef4501;
    assign array[34] = 32'h053775c0;
    assign array[35] = 32'h147d0004;
    assign array[36] = 32'hfc79239d;
    assign array[37] = 32'h441240a2;
    assign array[38] = 32'h80820131;
    assign array[39] = 32'hc2221151;
    assign array[40] = 32'hc026c406;
    assign array[41] = 32'h20000437;
    assign array[42] = 32'he9192a71;
    assign array[43] = 32'hfd6d2389;
    assign array[44] = 32'h44123f65;
    assign array[45] = 32'h448240a2;
    assign array[46] = 32'h20000337;
    assign array[47] = 32'h83020131;
    assign array[48] = 32'h225d8522;
    assign array[49] = 32'h00140493;
    assign array[50] = 32'h00080537;
    assign array[51] = 32'h84262b29;
    assign array[52] = 32'h1151bfe1;
    assign array[53] = 32'h2b9dc406;
    assign array[54] = 32'h40a23f41;
    assign array[55] = 32'h30000337;
    assign array[56] = 32'h83020131;
    assign array[57] = 32'hc8061131;
    assign array[58] = 32'hc426c622;
    assign array[59] = 32'h720000ef;
    assign array[60] = 32'hc00222b5;
    assign array[61] = 32'h04134782;
    assign array[62] = 32'h8b850400;
    assign array[63] = 32'ha03dc23e;
    assign array[64] = 32'h10000513;
    assign array[65] = 32'h21e521cd;
    assign array[66] = 32'h4792e50d;
    assign array[67] = 32'h0793c3a1;
    assign array[68] = 32'h85b30400;
    assign array[69] = 32'h8f854087;
    assign array[70] = 32'h00f5a5b3;
    assign array[71] = 32'h45014601;
    assign array[72] = 32'h00ef14fd;
    assign array[73] = 32'hfce96c00;
    assign array[74] = 32'hc81d147d;
    assign array[75] = 32'h04000493;
    assign array[76] = 32'h2a09bfc1;
    assign array[77] = 32'h4521d969;
    assign array[78] = 32'h4601297d;
    assign array[79] = 32'h45014581;
    assign array[80] = 32'h6a2000ef;
    assign array[81] = 32'hcd1d2201;
    assign array[82] = 32'ha0013f91;
    assign array[83] = 32'h04000793;
    assign array[84] = 32'h408785b3;
    assign array[85] = 32'ha5b38f85;
    assign array[86] = 32'hc59300f5;
    assign array[87] = 32'hbf7d0015;
    assign array[88] = 32'heb894792;
    assign array[89] = 32'h07854782;
    assign array[90] = 32'h4702c03e;
    assign array[91] = 32'h04e347c1;
    assign array[92] = 32'hb749fcf7;
    assign array[93] = 32'h00030537;
    assign array[94] = 32'h299521bd;
    assign array[95] = 32'h20d9d565;
    assign array[96] = 32'hbf55dd6d;
    assign array[97] = 32'hb7d137b9;
    assign array[98] = 32'h02054d63;
    assign array[99] = 32'hd3634799;
    assign array[100] = 32'h451900a7;
    assign array[101] = 32'h600007b7;
    assign array[102] = 32'h00b782a3;
    assign array[103] = 32'h06126585;
    assign array[104] = 32'h85930722;
    assign array[105] = 32'h7613f005;
    assign array[106] = 32'h8f6d0ff6;
    assign array[107] = 32'h8e498e59;
    assign array[108] = 32'h36b30642;
    assign array[109] = 32'h824100d0;
    assign array[110] = 32'h8e55068e;
    assign array[111] = 32'h00c79323;
    assign array[112] = 32'h45018082;
    assign array[113] = 32'h07b7bfc1;
    assign array[114] = 32'h43dc4000;
    assign array[115] = 32'h00a7d533;
    assign array[116] = 32'h80828905;
    assign array[117] = 32'h400007b7;
    assign array[118] = 32'h470543dc;
    assign array[119] = 32'h00a71533;
    assign array[120] = 32'h00e59763;
    assign array[121] = 32'h07378fc9;
    assign array[122] = 32'hc35c4000;
    assign array[123] = 32'h45138082;
    assign array[124] = 32'h8fe9fff5;
    assign array[125] = 32'h07b7bfcd;
    assign array[126] = 32'h439c4000;
    assign array[127] = 32'h00a7d533;
    assign array[128] = 32'h80828905;
    assign array[129] = 32'h95334785;
    assign array[130] = 32'hc59900a7;
    assign array[131] = 32'h40000737;
    assign array[132] = 32'h8d5d431c;
    assign array[133] = 32'h8082c308;
    assign array[134] = 32'h400007b7;
    assign array[135] = 32'h45134398;
    assign array[136] = 32'h8d79fff5;
    assign array[137] = 32'h8082c388;
    assign array[138] = 32'hc2221151;
    assign array[139] = 32'h842ac406;
    assign array[140] = 32'h459337d9;
    assign array[141] = 32'h85220015;
    assign array[142] = 32'h40a24412;
    assign array[143] = 32'h0ff5f593;
    assign array[144] = 32'hb7c90131;
    assign array[145] = 32'h500007b7;
    assign array[146] = 32'h0037c503;
    assign array[147] = 32'h80828905;
    assign array[148] = 32'h500007b7;
    assign array[149] = 32'h0027c503;
    assign array[150] = 32'h80828905;
    assign array[151] = 32'h500007b7;
    assign array[152] = 32'h81a34709;
    assign array[153] = 32'h808200e7;
    assign array[154] = 32'h4501e901;
    assign array[155] = 32'h45018082;
    assign array[156] = 32'h441240a2;
    assign array[157] = 32'h80820131;
    assign array[158] = 32'hc2221151;
    assign array[159] = 32'h842ac406;
    assign array[160] = 32'hd57537d1;
    assign array[161] = 32'h500007b7;
    assign array[162] = 32'h0017c783;
    assign array[163] = 32'h00f40023;
    assign array[164] = 32'h1151b7c5;
    assign array[165] = 32'hc406c222;
    assign array[166] = 32'h3f5d842a;
    assign array[167] = 32'h07b7c509;
    assign array[168] = 32'h80235000;
    assign array[169] = 32'h40a20087;
    assign array[170] = 32'h01314412;
    assign array[171] = 32'h11518082;
    assign array[172] = 32'hc026c222;
    assign array[173] = 32'h842ac406;
    assign array[174] = 32'h00b504b3;
    assign array[175] = 32'h00941763;
    assign array[176] = 32'h441240a2;
    assign array[177] = 32'h01314482;
    assign array[178] = 32'h85228082;
    assign array[179] = 32'hdd753f71;
    assign array[180] = 32'hb7ed0405;
    assign array[181] = 32'hc2221151;
    assign array[182] = 32'hc406c026;
    assign array[183] = 32'h04b3842a;
    assign array[184] = 32'h176300b5;
    assign array[185] = 32'h40a20094;
    assign array[186] = 32'h44824412;
    assign array[187] = 32'h80820131;
    assign array[188] = 32'h00044503;
    assign array[189] = 32'hdd6d3f79;
    assign array[190] = 32'hb7e50405;
    assign array[191] = 32'h600007b7;
    assign array[192] = 32'h0047c503;
    assign array[193] = 32'h3533897d;
    assign array[194] = 32'h808200a0;
    assign array[195] = 32'h600007b7;
    assign array[196] = 32'h0037c503;
    assign array[197] = 32'h3533897d;
    assign array[198] = 32'h808200a0;
    assign array[199] = 32'h600007b7;
    assign array[200] = 32'hf8000713;
    assign array[201] = 32'h00e78223;
    assign array[202] = 32'h07b78082;
    assign array[203] = 32'h07136000;
    assign array[204] = 32'h81a3f800;
    assign array[205] = 32'h808200e7;
    assign array[206] = 32'h4501e901;
    assign array[207] = 32'h45018082;
    assign array[208] = 32'h441240a2;
    assign array[209] = 32'h80820131;
    assign array[210] = 32'hc2221151;
    assign array[211] = 32'h842ac406;
    assign array[212] = 32'hd5753775;
    assign array[213] = 32'h600007b7;
    assign array[214] = 32'h0027c783;
    assign array[215] = 32'h00f40023;
    assign array[216] = 32'h1151b7c5;
    assign array[217] = 32'hc406c222;
    assign array[218] = 32'h374d842a;
    assign array[219] = 32'h07b7c509;
    assign array[220] = 32'h81236000;
    assign array[221] = 32'h40a20087;
    assign array[222] = 32'h01314412;
    assign array[223] = 32'h07b78082;
    assign array[224] = 32'hd5036000;
    assign array[225] = 32'h81050007;
    assign array[226] = 32'h80828905;
    assign array[227] = 32'h87936785;
    assign array[228] = 32'h059af007;
    assign array[229] = 32'h8d7d0522;
    assign array[230] = 32'h0ff5f593;
    assign array[231] = 32'he5938dc9;
    assign array[232] = 32'h07b70015;
    assign array[233] = 32'h90236000;
    assign array[234] = 32'h808200b7;
    assign array[235] = 32'h87936785;
    assign array[236] = 32'h059af007;
    assign array[237] = 32'h8d7d0522;
    assign array[238] = 32'h0ff5f593;
    assign array[239] = 32'he5938dc9;
    assign array[240] = 32'h07b70115;
    assign array[241] = 32'h90236000;
    assign array[242] = 32'h808200b7;
    assign array[243] = 32'h87936785;
    assign array[244] = 32'h059af007;
    assign array[245] = 32'h8d7d0522;
    assign array[246] = 32'h0ff5f593;
    assign array[247] = 32'he5938dc9;
    assign array[248] = 32'h07b70315;
    assign array[249] = 32'h90236000;
    assign array[250] = 32'h808200b7;
    assign array[251] = 32'h600007b7;
    assign array[252] = 32'h00079023;
    assign array[253] = 32'hc92d8082;
    assign array[254] = 32'hc8221121;
    assign array[255] = 32'hc626ca06;
    assign array[256] = 32'hc02ac232;
    assign array[257] = 32'hcd81842e;
    assign array[258] = 32'hfd7d3f9d;
    assign array[259] = 32'h600007b7;
    assign array[260] = 32'hf8000713;
    assign array[261] = 32'h00e78223;
    assign array[262] = 32'he7634481;
    assign array[263] = 32'h40d20084;
    assign array[264] = 32'h44b24442;
    assign array[265] = 32'h80820161;
    assign array[266] = 32'h409406b3;
    assign array[267] = 32'h73634741;
    assign array[268] = 32'h46c100d7;
    assign array[269] = 32'hf5134592;
    assign array[270] = 32'hc4360ff6;
    assign array[271] = 32'h46a23f81;
    assign array[272] = 32'h3f35c436;
    assign array[273] = 32'hfd6d46a2;
    assign array[274] = 32'h05374701;
    assign array[275] = 32'h47826000;
    assign array[276] = 32'h00254583;
    assign array[277] = 32'h00e48633;
    assign array[278] = 32'h0023963e;
    assign array[279] = 32'h070500b6;
    assign array[280] = 32'hfed717e3;
    assign array[281] = 32'hbf5594ba;
    assign array[282] = 32'hc92d8082;
    assign array[283] = 32'hc8221121;
    assign array[284] = 32'hc626ca06;
    assign array[285] = 32'hc02ac232;
    assign array[286] = 32'hcd81842e;
    assign array[287] = 32'hfd7d3709;
    assign array[288] = 32'h600007b7;
    assign array[289] = 32'hf8000713;
    assign array[290] = 32'h00e781a3;
    assign array[291] = 32'he7634481;
    assign array[292] = 32'h40d20084;
    assign array[293] = 32'h44b24442;
    assign array[294] = 32'h80820161;
    assign array[295] = 32'h40940733;
    assign array[296] = 32'hf36346c1;
    assign array[297] = 32'h474100e6;
    assign array[298] = 32'h05b74681;
    assign array[299] = 32'h47826000;
    assign array[300] = 32'h00d48633;
    assign array[301] = 32'h963e0685;
    assign array[302] = 32'h00064603;
    assign array[303] = 32'h00c58123;
    assign array[304] = 32'hfed717e3;
    assign array[305] = 32'h75134592;
    assign array[306] = 32'hc43a0ff7;
    assign array[307] = 32'h472235c5;
    assign array[308] = 32'h3575c43a;
    assign array[309] = 32'hfd6d4722;
    assign array[310] = 32'hbf5594ba;
    assign array[311] = 32'hcd358082;
    assign array[312] = 32'h0737cdad;
    assign array[313] = 32'h57836000;
    assign array[314] = 32'h8b890007;
    assign array[315] = 32'h0693ffed;
    assign array[316] = 32'h0223f800;
    assign array[317] = 32'h473d00d7;
    assign array[318] = 32'h06b77263;
    assign array[319] = 32'h00661713;
    assign array[320] = 32'h0ff77713;
    assign array[321] = 32'he7938fd9;
    assign array[322] = 32'h07370017;
    assign array[323] = 32'h10236000;
    assign array[324] = 32'h06b700f7;
    assign array[325] = 32'h47816000;
    assign array[326] = 32'h0046c703;
    assign array[327] = 32'h8b7d832e;
    assign array[328] = 32'h7363973e;
    assign array[329] = 32'h833a00b7;
    assign array[330] = 32'h0067fd63;
    assign array[331] = 32'h063397aa;
    assign array[332] = 32'hc7030065;
    assign array[333] = 32'h07850026;
    assign array[334] = 32'hfee78fa3;
    assign array[335] = 32'hfef61be3;
    assign array[336] = 32'hebe3879a;
    assign array[337] = 32'h0737fcb7;
    assign array[338] = 32'h57836000;
    assign array[339] = 32'h8b890007;
    assign array[340] = 32'h0793ffed;
    assign array[341] = 32'h0223f800;
    assign array[342] = 32'h808200f7;
    assign array[343] = 32'h00859793;
    assign array[344] = 32'h83c107c2;
    assign array[345] = 32'hc935bf61;
    assign array[346] = 32'h0737c9ad;
    assign array[347] = 32'h57836000;
    assign array[348] = 32'h8b890007;
    assign array[349] = 32'h0693ffed;
    assign array[350] = 32'h01a3f800;
    assign array[351] = 32'h473d00d7;
    assign array[352] = 32'h04b77e63;
    assign array[353] = 32'h00661713;
    assign array[354] = 32'h0ff77713;
    assign array[355] = 32'he7938fd9;
    assign array[356] = 32'h07370117;
    assign array[357] = 32'h10236000;
    assign array[358] = 32'h06b700f7;
    assign array[359] = 32'h47816000;
    assign array[360] = 32'h0036c703;
    assign array[361] = 32'h8b7d832e;
    assign array[362] = 32'h7363973e;
    assign array[363] = 32'h833a00b7;
    assign array[364] = 32'h0067fd63;
    assign array[365] = 32'h063397aa;
    assign array[366] = 32'hc7030065;
    assign array[367] = 32'h07850007;
    assign array[368] = 32'h00e68123;
    assign array[369] = 32'hfef61be3;
    assign array[370] = 32'hebe3879a;
    assign array[371] = 32'h0737fcb7;
    assign array[372] = 32'h57836000;
    assign array[373] = 32'h8b890007;
    assign array[374] = 32'h8082ffed;
    assign array[375] = 32'h00859793;
    assign array[376] = 32'h83c107c2;
    assign array[377] = 32'h07b7b745;
    assign array[378] = 32'hc3887000;
    assign array[379] = 32'h07b78082;
    assign array[380] = 32'h43887000;
    assign array[381] = 32'h07b78082;
    assign array[382] = 32'hc3887000;
    assign array[383] = 32'h70000737;
    assign array[384] = 32'hfffd431c;
    assign array[385] = 32'h07b78082;
    assign array[386] = 32'h8023f000;
    assign array[387] = 32'h80820007;
    assign array[388] = 32'hf00007b7;
    assign array[389] = 32'h80234705;
    assign array[390] = 32'h808200e7;
    assign array[391] = 32'hf00007b7;
    assign array[392] = 32'h8023471d;
    assign array[393] = 32'h808200e7;
    assign array[394] = 32'hf00007b7;
    assign array[395] = 32'h80234719;
    assign array[396] = 32'h808200e7;
    assign array[397] = 32'hf00007b7;
    assign array[398] = 32'h80234721;
    assign array[399] = 32'h808200e7;
    assign array[400] = 32'hf00007b7;
    assign array[401] = 32'h80234725;
    assign array[402] = 32'h808200e7;
    assign array[403] = 32'h4685470d;
    assign array[404] = 32'h05934611;
    assign array[405] = 32'h450d0bb0;
    assign array[406] = 32'h1141be05;
    assign array[407] = 32'hc422c606;
    assign array[408] = 32'h01051413;
    assign array[409] = 32'h31d13361;
    assign array[410] = 32'h45193955;
    assign array[411] = 32'h458139dd;
    assign array[412] = 32'h3b2d4505;
    assign array[413] = 32'h45293ba5;
    assign array[414] = 32'h05133fbd;
    assign array[415] = 32'h31d50d80;
    assign array[416] = 32'h01045513;
    assign array[417] = 32'h0ff57513;
    assign array[418] = 32'h450139e9;
    assign array[419] = 32'h450139d9;
    assign array[420] = 32'h458139c9;
    assign array[421] = 32'h3b194511;
    assign array[422] = 32'h45293b91;
    assign array[423] = 32'h45153fa9;
    assign array[424] = 32'h458131c9;
    assign array[425] = 32'h33194505;
    assign array[426] = 32'h45054581;
    assign array[427] = 32'h3b3d31c5;
    assign array[428] = 32'h00310513;
    assign array[429] = 32'h47833151;
    assign array[430] = 32'h8b850031;
    assign array[431] = 32'h40b2fff9;
    assign array[432] = 32'h01414422;
    assign array[433] = 32'h11118082;
    assign array[434] = 32'hca22cc06;
    assign array[435] = 32'hc22ec826;
    assign array[436] = 32'h0a058263;
    assign array[437] = 32'h0f6384b2;
    assign array[438] = 32'h14130806;
    assign array[439] = 32'hc0020085;
    assign array[440] = 32'h10000693;
    assign array[441] = 32'hf4638726;
    assign array[442] = 32'h07130096;
    assign array[443] = 32'hc43a1000;
    assign array[444] = 32'h392539f5;
    assign array[445] = 32'h45193125;
    assign array[446] = 32'h458131ad;
    assign array[447] = 32'h317d4505;
    assign array[448] = 32'h452931f5;
    assign array[449] = 32'h45093dcd;
    assign array[450] = 32'h551339a9;
    assign array[451] = 32'h75130104;
    assign array[452] = 32'h39810ff5;
    assign array[453] = 32'h00845513;
    assign array[454] = 32'h0ff57513;
    assign array[455] = 32'h75133199;
    assign array[456] = 32'h31810ff4;
    assign array[457] = 32'h45114581;
    assign array[458] = 32'h47223151;
    assign array[459] = 32'h46014792;
    assign array[460] = 32'h470285ba;
    assign array[461] = 32'h00e78533;
    assign array[462] = 32'h394d3b0d;
    assign array[463] = 32'h45294722;
    assign array[464] = 32'h3d55c43a;
    assign array[465] = 32'h39314515;
    assign array[466] = 32'h45054581;
    assign array[467] = 32'h45813185;
    assign array[468] = 32'h392d4505;
    assign array[469] = 32'h05133961;
    assign array[470] = 32'h3ef900f1;
    assign array[471] = 32'h00f14683;
    assign array[472] = 32'h8a854722;
    assign array[473] = 32'h4782fee9;
    assign array[474] = 32'h943a8c99;
    assign array[475] = 32'hc03e97ba;
    assign array[476] = 32'hf60498e3;
    assign array[477] = 32'h445240e2;
    assign array[478] = 32'h017144c2;
    assign array[479] = 32'hcdb98082;
    assign array[480] = 32'h1141ce31;
    assign array[481] = 32'hc032c606;
    assign array[482] = 32'hc226c422;
    assign array[483] = 32'h84ae842a;
    assign array[484] = 32'h3e6139b1;
    assign array[485] = 32'h05133661;
    assign array[486] = 32'h36e10bb0;
    assign array[487] = 32'h45054581;
    assign array[488] = 32'h55133131;
    assign array[489] = 32'h75130104;
    assign array[490] = 32'h3e650ff5;
    assign array[491] = 32'h00845513;
    assign array[492] = 32'h0ff57513;
    assign array[493] = 32'h7513367d;
    assign array[494] = 32'h36650ff4;
    assign array[495] = 32'h450d4585;
    assign array[496] = 32'h458536f5;
    assign array[497] = 32'h31194511;
    assign array[498] = 32'h85264782;
    assign array[499] = 32'h85be4605;
    assign array[500] = 32'h4422311d;
    assign array[501] = 32'h449240b2;
    assign array[502] = 32'hb9090141;
    assign array[503] = 32'h45018082;
    assign array[504] = 32'h1141bc19;
    assign array[505] = 32'h842ec422;
    assign array[506] = 32'h00154593;
    assign array[507] = 32'hc6064505;
    assign array[508] = 32'h3c09c032;
    assign array[509] = 32'h00144593;
    assign array[510] = 32'h34294509;
    assign array[511] = 32'h44224602;
    assign array[512] = 32'h459340b2;
    assign array[513] = 32'h450d0016;
    assign array[514] = 32'hbaed0141;
    assign array[515] = 32'h46011151;
    assign array[516] = 32'h45014581;
    assign array[517] = 32'h37f1c406;
    assign array[518] = 32'h45014581;
    assign array[519] = 32'h45853a65;
    assign array[520] = 32'h3a4d4505;
    assign array[521] = 32'h45094585;
    assign array[522] = 32'h40a23275;
    assign array[523] = 32'h450d4585;
    assign array[524] = 32'hb24d0131;
    assign array[525] = 32'h00000014;
    assign array[526] = 32'h00000000;
    assign array[527] = 32'h00527a01;
    assign array[528] = 32'h01017c01;
    assign array[529] = 32'h07020d1b;
    assign array[530] = 32'h00000001;
    assign array[531] = 32'h00000010;
    assign array[532] = 32'h0000001c;
    assign array[533] = 32'hfffff7ac;
    assign array[534] = 32'h00000016;
    assign array[535] = 32'h00000000;
