    assign array[0] = 32'h10001197;
    assign array[1] = 32'h80018193;
    assign array[2] = 32'h10000117;
    assign array[3] = 32'h1f810113;
    assign array[4] = 32'h11712015;
    assign array[5] = 32'h0040c022;
    assign array[6] = 32'hf00007b7;
    assign array[7] = 32'h00078023;
    assign array[8] = 32'h1171a001;
    assign array[9] = 32'h0040c022;
    assign array[10] = 32'hf00007b7;
    assign array[11] = 32'h80234705;
    assign array[12] = 32'ha00100e7;
    assign array[13] = 32'hc8061131;
    assign array[14] = 32'h0840c622;
    assign array[15] = 32'h600007b7;
    assign array[16] = 32'h30000713;
    assign array[17] = 32'h00e79323;
    assign array[18] = 32'h300007b7;
    assign array[19] = 32'h2823439c;
    assign array[20] = 32'h07b7fef4;
    assign array[21] = 32'h47096000;
    assign array[22] = 32'h00e78223;
    assign array[23] = 32'h600007b7;
    assign array[24] = 32'h8123470d;
    assign array[25] = 32'h07b700e7;
    assign array[26] = 32'h07136000;
    assign array[27] = 32'h90231050;
    assign array[28] = 32'h07b700e7;
    assign array[29] = 32'h81236000;
    assign array[30] = 32'h07b70007;
    assign array[31] = 32'h81236000;
    assign array[32] = 32'h07b70007;
    assign array[33] = 32'h81236000;
    assign array[34] = 32'h07b70007;
    assign array[35] = 32'h47156000;
    assign array[36] = 32'h00e79023;
    assign array[37] = 32'h600007b7;
    assign array[38] = 32'h82a34709;
    assign array[39] = 32'h07b700e7;
    assign array[40] = 32'h47056000;
    assign array[41] = 32'h00e79023;
    assign array[42] = 32'h600007b7;
    assign array[43] = 32'h00079023;
    assign array[44] = 32'hfe042623;
    assign array[45] = 32'h600007b7;
    assign array[46] = 32'h0037c783;
    assign array[47] = 32'h0ff7f793;
    assign array[48] = 32'h873e07e2;
    assign array[49] = 32'hfec42783;
    assign array[50] = 32'h8fd983a1;
    assign array[51] = 32'hfef42623;
    assign array[52] = 32'h600007b7;
    assign array[53] = 32'h0037c783;
    assign array[54] = 32'h0ff7f793;
    assign array[55] = 32'h873e07e2;
    assign array[56] = 32'hfec42783;
    assign array[57] = 32'h8fd983a1;
    assign array[58] = 32'hfef42623;
    assign array[59] = 32'h600007b7;
    assign array[60] = 32'h0037c783;
    assign array[61] = 32'h0ff7f793;
    assign array[62] = 32'h873e07e2;
    assign array[63] = 32'hfec42783;
    assign array[64] = 32'h8fd983a1;
    assign array[65] = 32'hfef42623;
    assign array[66] = 32'h600007b7;
    assign array[67] = 32'h0037c783;
    assign array[68] = 32'h0ff7f793;
    assign array[69] = 32'h873e07e2;
    assign array[70] = 32'hfec42783;
    assign array[71] = 32'h8fd983a1;
    assign array[72] = 32'hfef42623;
    assign array[73] = 32'h600007b7;
    assign array[74] = 32'h82a34709;
    assign array[75] = 32'h07b700e7;
    assign array[76] = 32'h27037000;
    assign array[77] = 32'hc398ff04;
    assign array[78] = 32'h700007b7;
    assign array[79] = 32'hfec42703;
    assign array[80] = 32'h2703c398;
    assign array[81] = 32'h2783ff04;
    assign array[82] = 32'h1463fec4;
    assign array[83] = 32'h35d100f7;
    assign array[84] = 32'h3dc1a011;
    assign array[85] = 32'h853e4781;
    assign array[86] = 32'h443240c2;
    assign array[87] = 32'h80820151;
    assign array[88] = 32'h00000014;
    assign array[89] = 32'h00000000;
    assign array[90] = 32'h00527a01;
    assign array[91] = 32'h01017c01;
    assign array[92] = 32'h07020d1b;
    assign array[93] = 32'h00000001;
    assign array[94] = 32'h00000010;
    assign array[95] = 32'h0000001c;
    assign array[96] = 32'hfffffe80;
    assign array[97] = 32'h00000012;
    assign array[98] = 32'h00000000;
